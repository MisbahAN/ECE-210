----------------------------------------------------------------------------------
-- Company: University of Alberta
-- Engineer: Behdad Goodarzy
-- 
-- Create Date: 09/06/2021 06:33:57 PM
-- Design Name: 
-- Module Name: tutorial - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity lab1 is
    Port ( sw : in STD_LOGIC_VECTOR (3 downto 0);
           led : out STD_LOGIC_VECTOR (1 downto 0)
           );
end lab1;

architecture Behavioral of lab1 is

begin
   
--
    
end Behavioral;
